module andm (inA, inB, out);
//1 bit and for (branch & zero)
input inA, inB;
output out;

assign out=inA&inB;

endmodule
